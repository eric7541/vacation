module top (
    input clk,
    input n_rst,
    input rxd,
    output txd
);

